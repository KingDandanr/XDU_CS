cpu5_inst : cpu5 PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
